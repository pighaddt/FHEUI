EX1                 ;第一行标题
VIN 1 0 AC 2V       ;独立电源说明，AC表示交流，2V表示幅值2V
R1 1 2 0.45K        ;电阻R1,阻值0.45k欧姆，连接节点1，2
R2 2 0 1K           ;电阻R2,1K欧姆，连接节点2，0
RI 3 0 1MEG         ;电阻RI，阻值1M欧姆(MEGA是10^3)，连接在节点3，0
R0 5 4 100          ;电阻R0,100欧姆，连接节点5，4
R3 3 4 500          ;电阻R3
R4 4 0 1K           ;电阻R4
C1 2 3 4U           ;电容C1，4微法，连接节点2，3
C2 2 4 4U           ;电容C2
E1 5 0 3 0 500K     ;电压控制电压源，系数A500k，输出端连接节点5，0，控制端连接节点3，0
.AC DEC 20 1 10K    ;DEC表示按数量级变化，20表示每一数量级取20个点，最后两个数表示起始频率和终止频率
                    *下面两条语句在ngspice没有用，*后面的也是注释，如果前面没有语句使用;做注释会报错
                    *.PLOT AC VM(4)     ;曲线打印语句，AC表示交流分析（正弦稳态分析），VM(4)表示节点4的电压 幅值
                    *.PROBE
.END                ;结束